`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:41:32 05/20/2023 
// Design Name: 
// Module Name:    MUX_16 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MUX_16(
    input [15:0] A0,
    input [15:0] A1,
    input sel,
    output [15:0] OUT
    );


endmodule
